`ifndef __ROB_SV__
`define __ROB_SV__
`include "ISA.svh"